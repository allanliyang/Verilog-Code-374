// T0: PCout, MARin, IncPC, Zin
// T1: Zlowout, PCin, MDMuxread, Mdatain, MDRin
// T2: MDRout, IRin
// T3: Grb, Rout, Yin
// T4: Cout, AND, Zin
// T5: Zlowout, Gra, Rin

// functionality
  // this tb performs addi R3, R4, 0x53
  // places result of (R4) && 0x53 in R3
`timescale 1ns/10ps
module datapath_tb_ANDI();
