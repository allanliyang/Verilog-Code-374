// T0: PCout, MARin, IncPC, Zin
// T1: Zlowout, PCin, MDMuxread, Mdatain, MDRin
// T2: MDRout, IRin
// T3: Grb, BAout, Yin
// T4: Cout, ADD, Zin
// T5: Zlowout, MARin
// T6: MDMuxread, Mdatain, MDRin
// T7: MDRout, Gra, Rin

// testbench for LD instruction
// NOTE: FIX TESTBENCH SETTINGS BEFORE RUNNING THIS

// functionality
	// this tb performs ld R2,0x95 and ld R0, 0x38(R2)
	
		
		
		
`timescale 1ns/10ps
module datapath_tb_LD();

endmodule
